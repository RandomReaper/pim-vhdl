-----------------------------------------------------------------------------
-- file			: tb.vhd 
--
-- brief		: Test bench
-- author(s)	: marc at pignat dot org
-- license		: The MIT License (MIT) (http://opensource.org/licenses/MIT)
--				  Copyright (c) 2015 Marc Pignat
-----------------------------------------------------------------------------

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
	
entity tb is
end tb;

architecture bhv of tb is
	signal reset			: std_ulogic;
	signal clock			: std_ulogic;
	signal adbus			: std_logic_vector(7 downto 0);
	signal txe_n			: std_ulogic;
	signal rxf_n			: std_ulogic;
	signal wr_n				: std_ulogic;
	signal rd_n				: std_ulogic;
	signal oe_n				: std_ulogic;
	signal siwu				: std_ulogic;
	signal suspend_n		: std_ulogic;
	signal reset_n			: std_ulogic;
	signal out_data_ack		: std_ulogic;
	signal counter			: unsigned(7 downto 0);
	signal out_data_write	: std_ulogic;
begin

reset_n <= not reset;

i_ft_if : entity work.ft245_sync_if
port map
(
	adbus			=> adbus,
	rxf_n			=> rxf_n,
	txe_n			=> txe_n,
	rd_n			=> rd_n,
	wr_n			=> wr_n,
	clkout			=> clock,
	oe_n			=> oe_n,
	siwu			=> siwu,
	reset_n			=> '0',
	suspend_n		=> suspend_n,
	
	reset			=> reset,
	in_data			=> open,
	in_data_read	=> '0',
	in_data_valid	=> open,
	
	out_data		=> std_ulogic_vector(counter),
	out_data_write	=> out_data_write,
	out_data_ack	=> out_data_ack
);

i_ft_sim : entity work.ft245_sync_sim
port map
(
	adbus		=> adbus,
	rxf_n		=> rxf_n,
	txe_n		=> txe_n,
	rd_n		=> rd_n,
	wr_n		=> wr_n,
	clkout		=> clock,
	oe_n		=> oe_n,
	siwu		=> siwu,
	reset_n		=> reset_n,
	suspend_n	=> suspend_n
);

i_reset : entity work.reset
port map
(
	reset	=> reset,
	clock	=> clock
);

counter_gen: process(reset, clock)
begin
	if reset = '1' then
		counter <= (others => '0');
		out_data_write <= '0';
	elsif rising_edge(clock) then
		out_data_write <= '0';
		if out_data_ack = '1' then
			counter <= counter + 1;
			out_data_write <= '1';
		end if;
	end if;
end process;

end bhv;